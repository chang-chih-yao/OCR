This is aaa.
!!!!
@@@
fksladjfl;dfjldfj
ieqru/cvj;gth]048510976
)~(@&*#(@&$_)!*(#@{%>?:"L{SDOGJKM