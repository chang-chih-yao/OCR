This is c.
skfjsalkfjlk
kdfja;slkdfjal;sf
kjasd;lfsakjdfl;aj
sjf;laskjdfl
132123165456411
1
32
132
132
1
231
3
46
54
89
74
[]
[
]\[
\[\
[\
(&*$#)(*@(*~&%)
19874-0`9240)!(*$&)(*$)?<?>S<?><
JLAK:SDFJLK:EJHRHIWHGOIDNND

